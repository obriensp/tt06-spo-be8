VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM16
  CLASS BLOCK ;
  FOREIGN RAM16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 111.320 BY 48.960 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 109.320 9.560 111.320 10.160 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 109.320 16.360 111.320 16.960 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 109.320 23.160 111.320 23.760 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 109.320 29.960 111.320 30.560 ;
    END
  END A0[3]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 109.320 36.760 111.320 37.360 ;
    END
  END CLK
  PIN Di0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 2.000 ;
    END
  END Di0[0]
  PIN Di0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 2.000 ;
    END
  END Di0[1]
  PIN Di0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 2.000 ;
    END
  END Di0[2]
  PIN Di0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 2.000 ;
    END
  END Di0[3]
  PIN Di0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 2.000 ;
    END
  END Di0[4]
  PIN Di0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 2.000 ;
    END
  END Di0[5]
  PIN Di0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 2.000 ;
    END
  END Di0[6]
  PIN Di0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 0.000 103.870 2.000 ;
    END
  END Di0[7]
  PIN Do0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 46.960 7.270 48.960 ;
    END
  END Do0[0]
  PIN Do0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 46.960 21.070 48.960 ;
    END
  END Do0[1]
  PIN Do0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 46.960 34.870 48.960 ;
    END
  END Do0[2]
  PIN Do0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 46.960 48.670 48.960 ;
    END
  END Do0[3]
  PIN Do0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 46.960 62.470 48.960 ;
    END
  END Do0[4]
  PIN Do0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 46.960 76.270 48.960 ;
    END
  END Do0[5]
  PIN Do0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 46.960 90.070 48.960 ;
    END
  END Do0[6]
  PIN Do0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 46.960 103.870 48.960 ;
    END
  END Do0[7]
  PIN EN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 109.320 2.760 111.320 3.360 ;
    END
  END EN0
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 92.320 -0.240 93.920 49.200 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 0.145 0.240 ;
    END
    PORT
      LAYER met1 ;
        RECT 111.175 -0.240 111.320 0.240 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 5.200 0.145 5.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 111.175 5.200 111.320 5.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 10.640 0.145 11.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 111.175 10.640 111.320 11.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 16.080 0.145 16.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 111.175 16.080 111.320 16.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 21.520 0.145 22.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 111.175 21.520 111.320 22.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 26.960 0.145 27.440 ;
    END
    PORT
      LAYER met1 ;
        RECT 111.175 26.960 111.320 27.440 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 32.400 0.145 32.880 ;
    END
    PORT
      LAYER met1 ;
        RECT 111.175 32.400 111.320 32.880 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 37.840 0.145 38.320 ;
    END
    PORT
      LAYER met1 ;
        RECT 111.175 37.840 111.320 38.320 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 43.280 0.145 43.760 ;
    END
    PORT
      LAYER met1 ;
        RECT 111.175 43.280 111.320 43.760 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 48.720 0.145 49.200 ;
    END
    PORT
      LAYER met1 ;
        RECT 111.175 48.720 111.320 49.200 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 15.520 -0.240 17.120 49.200 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 0.145 2.960 ;
    END
    PORT
      LAYER met1 ;
        RECT 111.175 2.480 111.320 2.960 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 7.920 0.145 8.400 ;
    END
    PORT
      LAYER met1 ;
        RECT 111.175 7.920 111.320 8.400 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 13.360 0.145 13.840 ;
    END
    PORT
      LAYER met1 ;
        RECT 111.175 13.360 111.320 13.840 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 18.800 0.145 19.280 ;
    END
    PORT
      LAYER met1 ;
        RECT 111.175 18.800 111.320 19.280 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 24.240 0.145 24.720 ;
    END
    PORT
      LAYER met1 ;
        RECT 111.175 24.240 111.320 24.720 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 29.680 0.145 30.160 ;
    END
    PORT
      LAYER met1 ;
        RECT 111.175 29.680 111.320 30.160 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 35.120 0.145 35.600 ;
    END
    PORT
      LAYER met1 ;
        RECT 111.175 35.120 111.320 35.600 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 40.560 0.145 41.040 ;
    END
    PORT
      LAYER met1 ;
        RECT 111.175 40.560 111.320 41.040 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 46.000 0.145 46.480 ;
    END
    PORT
      LAYER met1 ;
        RECT 111.175 46.000 111.320 46.480 ;
    END
  END VPWR
  PIN WE0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 109.320 43.560 111.320 44.160 ;
    END
  END WE0
  OBS
      LAYER pwell ;
        RECT 0.605 48.855 0.775 49.045 ;
        RECT 3.365 48.855 3.535 49.045 ;
        RECT 6.125 48.855 6.295 49.045 ;
        RECT 13.485 48.895 13.655 49.045 ;
        RECT 14.865 48.855 15.035 49.045 ;
        RECT 22.225 48.895 22.395 49.045 ;
        RECT 23.605 48.855 23.775 49.045 ;
        RECT 30.965 48.895 31.135 49.045 ;
        RECT 32.345 48.855 32.515 49.045 ;
        RECT 39.705 48.895 39.875 49.045 ;
        RECT 41.085 48.855 41.255 49.045 ;
        RECT 48.445 48.895 48.615 49.045 ;
        RECT 49.825 48.855 49.995 49.045 ;
        RECT 57.185 48.895 57.355 49.045 ;
        RECT 58.565 48.855 58.735 49.045 ;
        RECT 65.925 48.895 66.095 49.045 ;
        RECT 67.305 48.855 67.475 49.045 ;
        RECT 74.665 48.895 74.835 49.045 ;
        RECT 76.045 48.855 76.215 49.045 ;
        RECT 81.565 48.855 81.735 49.045 ;
        RECT 87.545 48.855 87.715 49.045 ;
        RECT 93.065 48.855 93.235 49.045 ;
        RECT 99.045 48.855 99.215 49.045 ;
        RECT 104.565 48.855 104.735 49.045 ;
        RECT 108.705 48.855 108.875 49.045 ;
      LAYER nwell ;
        RECT -0.190 44.825 111.510 47.655 ;
        RECT -0.190 42.165 82.415 42.215 ;
        RECT 84.040 42.165 111.510 42.215 ;
        RECT -0.190 39.435 111.510 42.165 ;
        RECT -0.190 39.385 81.955 39.435 ;
        RECT 83.580 39.385 111.510 39.435 ;
        RECT -0.190 36.725 82.415 36.775 ;
        RECT 84.040 36.725 111.510 36.775 ;
        RECT -0.190 33.995 111.510 36.725 ;
        RECT -0.190 33.945 81.955 33.995 ;
        RECT 83.580 33.945 111.510 33.995 ;
        RECT -0.190 31.285 82.415 31.335 ;
        RECT 84.040 31.285 111.510 31.335 ;
        RECT -0.190 28.555 111.510 31.285 ;
        RECT -0.190 28.505 81.955 28.555 ;
        RECT 83.580 28.505 111.510 28.555 ;
        RECT -0.190 25.845 82.415 25.895 ;
        RECT 84.040 25.845 111.510 25.895 ;
        RECT -0.190 23.115 111.510 25.845 ;
        RECT -0.190 23.065 81.955 23.115 ;
        RECT 83.580 23.065 111.510 23.115 ;
        RECT -0.190 20.405 82.415 20.455 ;
        RECT 84.040 20.405 111.510 20.455 ;
        RECT -0.190 17.675 111.510 20.405 ;
        RECT -0.190 17.625 81.955 17.675 ;
        RECT 83.580 17.625 111.510 17.675 ;
        RECT -0.190 14.965 82.415 15.015 ;
        RECT 84.040 14.965 111.510 15.015 ;
        RECT -0.190 12.235 111.510 14.965 ;
        RECT -0.190 12.185 81.955 12.235 ;
        RECT 83.580 12.185 111.510 12.235 ;
        RECT -0.190 9.525 82.415 9.575 ;
        RECT 84.040 9.525 111.510 9.575 ;
        RECT -0.190 6.795 111.510 9.525 ;
        RECT -0.190 6.745 81.955 6.795 ;
        RECT 83.580 6.745 111.510 6.795 ;
        RECT -0.190 4.085 82.415 4.135 ;
        RECT 84.040 4.085 111.510 4.135 ;
        RECT -0.190 1.355 111.510 4.085 ;
        RECT -0.190 1.305 81.955 1.355 ;
        RECT 83.580 1.305 111.510 1.355 ;
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.105 ;
        RECT 5.670 -0.085 5.840 0.105 ;
        RECT 10.265 -0.085 10.435 0.105 ;
        RECT 15.790 -0.085 15.960 0.105 ;
        RECT 20.385 -0.085 20.555 0.105 ;
        RECT 25.910 -0.085 26.080 0.105 ;
        RECT 30.505 -0.085 30.675 0.105 ;
        RECT 36.030 -0.085 36.200 0.105 ;
        RECT 40.625 -0.085 40.795 0.105 ;
        RECT 46.150 -0.085 46.320 0.105 ;
        RECT 50.745 -0.085 50.915 0.105 ;
        RECT 56.270 -0.085 56.440 0.105 ;
        RECT 60.865 -0.085 61.035 0.105 ;
        RECT 66.390 -0.085 66.560 0.105 ;
        RECT 70.985 -0.085 71.155 0.105 ;
        RECT 76.510 -0.085 76.680 0.105 ;
        RECT 81.110 -0.085 81.280 0.105 ;
        RECT 87.545 -0.085 87.715 0.085 ;
        RECT 89.845 -0.085 90.015 0.065 ;
        RECT 90.765 -0.085 90.935 0.085 ;
        RECT 92.145 -0.085 92.315 0.085 ;
        RECT 93.985 -0.085 94.155 0.105 ;
        RECT 96.745 -0.085 96.915 0.105 ;
        RECT 99.045 -0.085 99.215 0.105 ;
        RECT 100.885 -0.085 101.055 0.105 ;
        RECT 106.405 -0.085 106.575 0.105 ;
        RECT 108.245 -0.085 108.415 0.105 ;
        RECT 110.555 -0.050 110.715 0.060 ;
      LAYER li1 ;
        RECT 0.000 48.875 111.320 49.045 ;
      LAYER li1 ;
        RECT 0.000 0.085 111.320 48.875 ;
      LAYER li1 ;
        RECT 0.000 -0.085 111.320 0.085 ;
      LAYER met1 ;
        RECT 0.145 48.875 111.175 49.200 ;
        RECT 0.425 48.440 110.895 48.875 ;
        RECT 0.085 46.760 111.175 48.440 ;
        RECT 0.425 45.720 110.895 46.760 ;
        RECT 0.085 44.040 111.175 45.720 ;
        RECT 0.425 43.000 110.895 44.040 ;
        RECT 0.085 41.320 111.175 43.000 ;
        RECT 0.425 40.280 110.895 41.320 ;
        RECT 0.085 38.600 111.175 40.280 ;
        RECT 0.425 37.560 110.895 38.600 ;
        RECT 0.085 35.880 111.175 37.560 ;
        RECT 0.425 34.840 110.895 35.880 ;
        RECT 0.085 33.160 111.175 34.840 ;
        RECT 0.425 32.120 110.895 33.160 ;
        RECT 0.085 30.440 111.175 32.120 ;
        RECT 0.425 29.400 110.895 30.440 ;
        RECT 0.085 27.720 111.175 29.400 ;
        RECT 0.425 26.680 110.895 27.720 ;
        RECT 0.085 25.000 111.175 26.680 ;
        RECT 0.425 23.960 110.895 25.000 ;
        RECT 0.085 22.280 111.175 23.960 ;
        RECT 0.425 21.240 110.895 22.280 ;
        RECT 0.085 19.560 111.175 21.240 ;
        RECT 0.425 18.520 110.895 19.560 ;
        RECT 0.085 16.840 111.175 18.520 ;
        RECT 0.425 15.800 110.895 16.840 ;
        RECT 0.085 14.120 111.175 15.800 ;
        RECT 0.425 13.080 110.895 14.120 ;
        RECT 0.085 11.400 111.175 13.080 ;
        RECT 0.425 10.360 110.895 11.400 ;
        RECT 0.085 8.680 111.175 10.360 ;
        RECT 0.425 7.640 110.895 8.680 ;
        RECT 0.085 5.960 111.175 7.640 ;
        RECT 0.425 4.920 110.895 5.960 ;
        RECT 0.085 3.240 111.175 4.920 ;
        RECT 0.425 2.200 110.895 3.240 ;
        RECT 0.085 0.520 111.175 2.200 ;
        RECT 0.425 0.085 110.895 0.520 ;
        RECT 0.145 -0.240 111.175 0.085 ;
      LAYER met2 ;
        RECT 92.350 48.960 93.890 49.145 ;
        RECT 1.940 46.680 6.710 48.960 ;
        RECT 7.550 46.680 20.510 48.960 ;
        RECT 21.350 46.680 34.310 48.960 ;
        RECT 35.150 46.680 48.110 48.960 ;
        RECT 48.950 46.680 61.910 48.960 ;
        RECT 62.750 46.680 75.710 48.960 ;
        RECT 76.550 46.680 89.510 48.960 ;
        RECT 90.350 46.680 103.310 48.960 ;
        RECT 104.150 46.680 110.760 48.960 ;
        RECT 1.940 2.280 110.760 46.680 ;
        RECT 1.940 0.000 6.710 2.280 ;
        RECT 7.550 0.000 20.510 2.280 ;
        RECT 21.350 0.000 34.310 2.280 ;
        RECT 35.150 0.000 48.110 2.280 ;
        RECT 48.950 0.000 61.910 2.280 ;
        RECT 62.750 0.000 75.710 2.280 ;
        RECT 76.550 0.000 89.510 2.280 ;
        RECT 90.350 0.000 103.310 2.280 ;
        RECT 104.150 0.000 110.760 2.280 ;
        RECT 92.350 -0.185 93.890 0.000 ;
      LAYER met3 ;
        RECT 92.330 48.960 93.910 49.125 ;
        RECT 13.865 44.560 109.320 48.960 ;
        RECT 13.865 43.160 108.920 44.560 ;
        RECT 13.865 37.760 109.320 43.160 ;
        RECT 13.865 36.360 108.920 37.760 ;
        RECT 13.865 30.960 109.320 36.360 ;
        RECT 13.865 29.560 108.920 30.960 ;
        RECT 13.865 24.160 109.320 29.560 ;
        RECT 13.865 22.760 108.920 24.160 ;
        RECT 13.865 17.360 109.320 22.760 ;
        RECT 13.865 15.960 108.920 17.360 ;
        RECT 13.865 10.560 109.320 15.960 ;
        RECT 13.865 9.160 108.920 10.560 ;
        RECT 13.865 3.760 109.320 9.160 ;
        RECT 13.865 2.360 108.920 3.760 ;
        RECT 13.865 0.000 109.320 2.360 ;
        RECT 92.330 -0.165 93.910 0.000 ;
  END
END RAM16
END LIBRARY

